module led(clk,row,col,w);           
input clk;                    
output [15:0] row;               
output [3:0] col;                 
reg [3:0] col;
reg [15:0] row;
input [2:0]w;

always @(posedge clk)
	begin
	case(w)
	3'b000:begin
	case(col)                                       
	4'b0000:row<=16'b0000000000000000;
	4'b0001:row<=16'b0000000000000000;
	4'b0010:row<=16'b0000000000000000;
	4'b0011:row<=16'b0000000000000000;
	4'b0100:row<=16'b0000000000000000;
	4'b0101:row<=16'b0000000000000000;
	4'b0110:row<=16'b0000000000000000;
	4'b0111:row<=16'b0000000000000000;
	4'b1000:row<=16'b0000000000000000;
	4'b1001:row<=16'b0000000000000000;
	4'b1010:row<=16'b0000000000000000;
	4'b1011:row<=16'b0000000000000000;
	4'b1100:row<=16'b0000000000000000;
	4'b1101:row<=16'b0000000000000000;
	4'b1110:row<=16'b0000000000000000;
	4'b1111:row<=16'b0000000000000000;
	endcase
	end
	
	3'b001:begin
	case(col)                                       
	4'b0000:row<=16'b0000000000000000;
	4'b0001:row<=16'b0000000000000000;
	4'b0010:row<=16'b0000000000000000;
	4'b0011:row<=16'b0000000000000000;
	4'b0100:row<=16'b0000000000000000;
	4'b0101:row<=16'b0000000000000000;
	4'b0110:row<=16'b0000000000000000;
	4'b0111:row<=16'b1111111111111111;
	4'b1000:row<=16'b0000000000000000;
	4'b1001:row<=16'b0000000000000000;
	4'b1010:row<=16'b0000000000000000;
	4'b1011:row<=16'b0000000000000000;
	4'b1100:row<=16'b0000000000000000;
	4'b1101:row<=16'b0000000000000000;
	4'b1110:row<=16'b0000000000000000;
	4'b1111:row<=16'b0000000000000000;
	endcase
	end
	
	3'b010:begin
	case(col)                                       
	4'b0000:row<=16'b0000000000000000;
	4'b0001:row<=16'b0000000000000000;
	4'b0010:row<=16'b0000000000000000;
	4'b0011:row<=16'b0000000000000000;
	4'b0100:row<=16'b0011111111111100;
	4'b0101:row<=16'b0000000000000000;
	4'b0110:row<=16'b0000000000000000;
	4'b0111:row<=16'b0000000000000000;
	4'b1000:row<=16'b0000000000000000;
	4'b1001:row<=16'b0000000000000000;
	4'b1010:row<=16'b1111111111111111;
	4'b1011:row<=16'b0000000000000000;
	4'b1100:row<=16'b0000000000000000;
	4'b1101:row<=16'b0000000000000000;
	4'b1110:row<=16'b0000000000000000;
	4'b1111:row<=16'b0000000000000000;
	endcase
	end
	
	3'b011:begin
	case(col)                                       
	4'b0000:row<=16'b0000000000000000;
	4'b0001:row<=16'b0000000000000000;
	4'b0010:row<=16'b0000000000000000;
	4'b0011:row<=16'b0011111111111100;
	4'b0100:row<=16'b0000000000000000;
	4'b0101:row<=16'b0000000000000000;
	4'b0110:row<=16'b0000111111110000;
	4'b0111:row<=16'b0000000000000000;
	4'b1000:row<=16'b0000000000000000;
	4'b1001:row<=16'b0000000000000000;
	4'b1010:row<=16'b1111111111111111;
	4'b1011:row<=16'b0000000000000000;
	4'b1100:row<=16'b0000000000000000;
	4'b1101:row<=16'b0000000000000000;
	4'b1110:row<=16'b0000000000000000;
	4'b1111:row<=16'b0000000000000000;
	endcase
	end
	
	3'b100:begin
	case(col)                                       
	4'b0000:row<=16'b0000000000000000;
	4'b0001:row<=16'b0000000000000000;
	4'b0010:row<=16'b0000000000000000;
	4'b0011:row<=16'b1111111111111111;
	4'b0100:row<=16'b1000010000100001;
	4'b0101:row<=16'b1000010000100001;
	4'b0110:row<=16'b1000010000100001;
	4'b0111:row<=16'b1111110000111111;
	4'b1000:row<=16'b1000000000000001;
	4'b1001:row<=16'b1000000000000001;
	4'b1010:row<=16'b1000000000000001;
	4'b1011:row<=16'b1111111111111111;
	4'b1100:row<=16'b0000000000000000;
	4'b1101:row<=16'b0000000000000000;
	4'b1110:row<=16'b0000000000000000;
	4'b1111:row<=16'b0000000000000000;
	endcase
	end
	
	default:begin 
	case(col)                                       
	4'b0000:row<=16'b0000000000000000;
	4'b0001:row<=16'b0000000000000000;
	4'b0010:row<=16'b0000000000000000;
	4'b0011:row<=16'b0000000000000000;
	4'b0100:row<=16'b0000000000000000;
	4'b0101:row<=16'b0000000000000000;
	4'b0110:row<=16'b0000000000000000;
	4'b0111:row<=16'b0000000000000000;
	4'b1000:row<=16'b0000000000000000;
	4'b1001:row<=16'b0000000000000000;
	4'b1010:row<=16'b0000000000000000;
	4'b1011:row<=16'b0000000000000000;
	4'b1100:row<=16'b0000000000000000;
	4'b1101:row<=16'b0000000000000000;
	4'b1110:row<=16'b0000000000000000;
	4'b1111:row<=16'b0000000000000000;
	endcase		
	end
	endcase
	end
	
	always@(posedge clk)
	begin
	case(col)                                              
	4'b0000:col<=4'b0001;
	4'b0001:col<=4'b0010;
	4'b0010:col<=4'b0011;
	4'b0011:col<=4'b0100;
	4'b0100:col<=4'b0101;
	4'b0101:col<=4'b0110;
	4'b0110:col<=4'b0111;
	4'b0111:col<=4'b1000;
	4'b1000:col<=4'b1001;
	4'b1001:col<=4'b1010;
	4'b1010:col<=4'b1011;
	4'b1011:col<=4'b1100;
	4'b1100:col<=4'b1101;
	4'b1101:col<=4'b1110;
	4'b1110:col<=4'b1111;
	4'b1111:col<=4'b0000;
	default:col<=4'b0000;
	endcase
	end
	
	endmodule
	
	