module led(clk,row,col);           
input clk;                    
output [15:0] row;               
output [3:0] col;                 
reg [3:0] col;
reg [15:0] row;
always @(posedge clk)
	begin
	case(col)                                       
	4'b0000:row<=16'b0000000000000000;
	4'b0001:row<=16'b0000000000000000;
	4'b0010:row<=16'b0000000000000000;
	4'b0011:row<=16'b0000000000000000;
	4'b0100:row<=16'b0000000000000000;
	4'b0101:row<=16'b0000000000000000;
	4'b0110:row<=16'b0000000000000000;
	4'b0111:row<=16'b0000000000000000;
	4'b1000:row<=16'b0000000000000000;
	4'b1001:row<=16'b0000000000000000;
	4'b1010:row<=16'b0000000000000000;
	4'b1011:row<=16'b0000000000000000;
	4'b1100:row<=16'b0000000000000000;
	4'b1101:row<=16'b0000000000000000;
	4'b1110:row<=16'b0000000000000000;
	4'b1111:row<=16'b0000000000000000;
	endcase
	end
	
	always@(posedge clk)
	begin
	case(col)                                              
	4'b0000:col<=4'b0001;
	4'b0001:col<=4'b0010;
	4'b0010:col<=4'b0011;
	4'b0011:col<=4'b0100;
	4'b0100:col<=4'b0101;
	4'b0101:col<=4'b0110;
	4'b0110:col<=4'b0111;
	4'b0111:col<=4'b1000;
	4'b1000:col<=4'b1001;
	4'b1001:col<=4'b1010;
	4'b1010:col<=4'b1011;
	4'b1011:col<=4'b1100;
	4'b1100:col<=4'b1101;
	4'b1101:col<=4'b1110;
	4'b1110:col<=4'b1111;
	4'b1111:col<=4'b0000;
	default:col<=4'b0000;
	endcase
	end
	
	endmodule
	
	