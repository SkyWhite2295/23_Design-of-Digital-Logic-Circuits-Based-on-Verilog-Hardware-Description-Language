module show_score(p1_s,p2_s,p3_s,p4_s,d0,d1,d2,d3,d4,d5,d6,d7,h);
wire h;
assign h = 1'b0;
input [3:0]p1_s,p2_s,p3_s,p4_s;
output h;
output [3:0]d0,d1,d2,d3,d4,d5,d6,d7;
reg [3:0]d0,d1,d2,d3,d4,d5,d6,d7;

always @ (p1_s)
begin
case(p1_s)
4'b0000:{d7,d6}=8'b00000000;
4'b0001:{d7,d6}=8'b00000001;
4'b0010:{d7,d6}=8'b00000010;
4'b0011:{d7,d6}=8'b00000011;
4'b0100:{d7,d6}=8'b00000100;
4'b0101:{d7,d6}=8'b00000101;
4'b0110:{d7,d6}=8'b00000110;
4'b0111:{d7,d6}=8'b00000111;
4'b1000:{d7,d6}=8'b00001000;
4'b1001:{d7,d6}=8'b00001001;
4'b1010:{d7,d6}=8'b00010000;
4'b1011:{d7,d6}=8'b00010001;
4'b1100:{d7,d6}=8'b00010010;
4'b1101:{d7,d6}=8'b00010011;
4'b1110:{d7,d6}=8'b00010100;
4'b1111:{d7,d6}=8'b00010101;
default:{d7,d6}=8'b00000000;
endcase
end

always @ (p2_s)
begin
case(p2_s)
4'b0000:{d5,d4}=8'b00000000;
4'b0001:{d5,d4}=8'b00000001;
4'b0010:{d5,d4}=8'b00000010;
4'b0011:{d5,d4}=8'b00000011;
4'b0100:{d5,d4}=8'b00000100;
4'b0101:{d5,d4}=8'b00000101;
4'b0110:{d5,d4}=8'b00000110;
4'b0111:{d5,d4}=8'b00000111;
4'b1000:{d5,d4}=8'b00001000;
4'b1001:{d5,d4}=8'b00001001;
4'b1010:{d5,d4}=8'b00010000;
4'b1011:{d5,d4}=8'b00010001;
4'b1100:{d5,d4}=8'b00010010;
4'b1101:{d5,d4}=8'b00010011;
4'b1110:{d5,d4}=8'b00010100;
4'b1111:{d5,d4}=8'b00010101;
default:{d5,d4}=8'b00000000;
endcase
end

always @ (p3_s)
begin
case(p3_s)
4'b0000:{d3,d2}=8'b00000000;
4'b0001:{d3,d2}=8'b00000001;
4'b0010:{d3,d2}=8'b00000010;
4'b0011:{d3,d2}=8'b00000011;
4'b0100:{d3,d2}=8'b00000100;
4'b0101:{d3,d2}=8'b00000101;
4'b0110:{d3,d2}=8'b00000110;
4'b0111:{d3,d2}=8'b00000111;
4'b1000:{d3,d2}=8'b00001000;
4'b1001:{d3,d2}=8'b00001001;
4'b1010:{d3,d2}=8'b00010000;
4'b1011:{d3,d2}=8'b00010001;
4'b1100:{d3,d2}=8'b00010010;
4'b1101:{d3,d2}=8'b00010011;
4'b1110:{d3,d2}=8'b00010100;
4'b1111:{d3,d2}=8'b00010101;
default:{d3,d2}=8'b00000000;
endcase
end

always @ (p4_s)
begin
case(p4_s)
4'b0000:{d1,d0}=8'b00000000;
4'b0001:{d1,d0}=8'b00000001;
4'b0010:{d1,d0}=8'b00000010;
4'b0011:{d1,d0}=8'b00000011;
4'b0100:{d1,d0}=8'b00000100;
4'b0101:{d1,d0}=8'b00000101;
4'b0110:{d1,d0}=8'b00000110;
4'b0111:{d1,d0}=8'b00000111;
4'b1000:{d1,d0}=8'b00001000;
4'b1001:{d1,d0}=8'b00001001;
4'b1010:{d1,d0}=8'b00010000;
4'b1011:{d1,d0}=8'b00010001;
4'b1100:{d1,d0}=8'b00010010;
4'b1101:{d1,d0}=8'b00010011;
4'b1110:{d1,d0}=8'b00010100;
4'b1111:{d1,d0}=8'b00010101;
default:{d1,d0}=8'b00000000;
endcase
end

endmodule
